200
33 4 12 23 108 r 50 45 42 34 h 23 T 35 H 46 T 50 H 52 B
50 34 9 42 20 r h 39 B 44 B
47 45 37 52 69 r h 0 B 32 B
30 0 56 5 62 r h 8 B 20 B
0 3 1 10 3 5 1 4 5 7 3 10 2 11 0 3 3 8 0 2 0 6 1 8 4 12 1 5 4 11 2 4 4 6 2 9 2 9 
15
